`timescale 1ns / 1ps

////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer:
//
// Create Date:   21:49:27 12/09/2017
// Design Name:   file
// Module Name:   E:/ISEproject/fileIOtest/IOtest.v
// Project Name:  fileIOtest
// Target Device:  
// Tool versions:  
// Description: 
//
// Verilog Test Fixture created by ISE for module: file
//
// Dependencies:
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
////////////////////////////////////////////////////////////////////////////////

module IOtest;

	// Outputs
	wire [31:0] out;

	// Instantiate the Unit Under Test (UUT)
	file uut (
		.out(out)
	);

	initial begin
		// Initialize Inputs

		// Wait 100 ns for global reset to finish
		
        
		// Add stimulus here

	end
      
endmodule

